// VGA protocol constants for 800x600 resolution
`define VGA_WIDTH  800
`define VGA_HEIGHT 600
`define VGA_HLIMIT 1056
`define VGA_VLIMIT 628
`define VGA_HSYNC_PULSE_START 840
`define VGA_HSYNC_PULSE_END   968
`define VGA_VSYNC_PULSE_START 601
`define VGA_VSYNC_PULSE_END   605

`define IMAGEN_PIXELS 15000
`define IMAGE_WIDTH 150
`define IMAGE_HEIGHT 100

`define POSITION_H 290
`define POSITION_V 200

`define RED 8'he0;
`define GREEN 8'h1c
`define BLUE 8'h3
`define BLANK 8'hff
`define BLACK 8'h00

`define COLOR_BITS 8
